`timescale 1ns / 1ps

// �Ĵ����ļ���Ҫ���logisim�ϵ���ȫ��ͬ
module RegFile();
endmodule
