`timescale 1ns / 1ps
// ��������������뱣֤��ȷ
module AluController(

    );
endmodule
