`timescale 1ns / 1ps

// �����������������logisim�ϵ���ͬ
module ALU();
endmodule
