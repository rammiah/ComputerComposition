`timescale 1ns / 1ps
// �޷��űȽ�������logisim��ͬ
module UCompare();
endmodule
