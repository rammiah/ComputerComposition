`timescale 1ns / 1ps
// ��·ѡ������ѡ���ź�Ϊ1λ�ģ�����2������
module MUX2();
endmodule
