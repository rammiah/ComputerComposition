`timescale 1ns / 1ps
// �����űȽ�������logisim��ͬ
module Compare(

    );
endmodule
