`timescale 1ns / 1ps
// �����ź����ɣ�������ȷ
module ControlSignal(

    );
endmodule
