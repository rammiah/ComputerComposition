`timescale 1ns / 1ps

module LRightShifter(

    );
endmodule
