`timescale 1ns / 1ps
// ��չ�ź����ɣ������Լ�д�Լ���
module ExtendSignal();
endmodule
