`timescale 1ns / 1ps
// ʵ��mips-ram��Ҫ���logisim��ȫ��ͬ��
// ʹ��˵��д���ĵ���,RAM���Բ�����
module RAM();
endmodule
