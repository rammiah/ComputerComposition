`timescale 1ns / 1ps
// ������չ
module SignedExt(

    );
endmodule
