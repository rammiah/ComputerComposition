`timescale 1ns / 1ps
// ������������ʵ��logisim��ԭ�ȸ��Ľӿڣ�Ԥ��4���������չָ�c1, c2, m, b
module Controller();
endmodule
