`timescale 1ns / 1ps
// ��������ʱ�������ؼ�����һ��rst��λ,ʵ��logisim��
// �еļ��������ɣ�����Ҫ���� -1
module Counter();
endmodule
