`timescale 1ns / 1ps
// ��·ѡ����������ѡ���ź�Ϊ2λ
module MUX4();

endmodule
