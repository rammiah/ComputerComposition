`timescale 1ns / 1ps
// �޷�����չ
module UnsignedExt(

    );
endmodule
