`timescale 1ns / 1ps
// ʵ��PC�Ĵ���
module PC(

    );
endmodule
