`timescale 1ns / 1ps
// �����Լ�����Լ��ģ������Լ�����չָ�����
module CPU();
// �������

endmodule
